-------------------------------------------------------------------------
-- Sullivan Hart
-------------------------------------------------------------------------
-- decoder5bit.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of a 5 bit to 32 bit decoder
-------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY decoder5bit IS
	PORT (
		i_In : IN STD_LOGIC_VECTOR(4 DOWNTO 0); -- Data value input
		i_En : IN STD_LOGIC;
		o_Out : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)); -- Data value output

END decoder5bit;

ARCHITECTURE mixed OF decoder5bit IS

	COMPONENT mux2t1_N
		PORT (
			i_S : IN STD_LOGIC;
			i_D0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			i_D1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			o_O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
	END COMPONENT;

	SIGNAL decoderOut : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN

	WITH i_In SELECT
		decoderOut <=

		"00000000000000000000000000000001" WHEN "00000",
		"00000000000000000000000000000010" WHEN "00001",
		"00000000000000000000000000000100" WHEN "00010",
		"00000000000000000000000000001000" WHEN "00011",
		"00000000000000000000000000010000" WHEN "00100",
		"00000000000000000000000000100000" WHEN "00101",
		"00000000000000000000000001000000" WHEN "00110",
		"00000000000000000000000010000000" WHEN "00111",
		"00000000000000000000000100000000" WHEN "01000",
		"00000000000000000000001000000000" WHEN "01001",
		"00000000000000000000010000000000" WHEN "01010",
		"00000000000000000000100000000000" WHEN "01011",
		"00000000000000000001000000000000" WHEN "01100",
		"00000000000000000010000000000000" WHEN "01101",
		"00000000000000000100000000000000" WHEN "01110",
		"00000000000000001000000000000000" WHEN "01111",
		"00000000000000010000000000000000" WHEN "10000",
		"00000000000000100000000000000000" WHEN "10001",
		"00000000000001000000000000000000" WHEN "10010",
		"00000000000010000000000000000000" WHEN "10011",
		"00000000000100000000000000000000" WHEN "10100",
		"00000000001000000000000000000000" WHEN "10101",
		"00000000010000000000000000000000" WHEN "10110",
		"00000000100000000000000000000000" WHEN "10111",
		"00000001000000000000000000000000" WHEN "11000",
		"00000010000000000000000000000000" WHEN "11001",
		"00000100000000000000000000000000" WHEN "11010",
		"00001000000000000000000000000000" WHEN "11011",
		"00010000000000000000000000000000" WHEN "11100",
		"00100000000000000000000000000000" WHEN "11101",
		"01000000000000000000000000000000" WHEN "11110",
		"10000000000000000000000000000000" WHEN "11111",
		"00000000000000000000000000000000" WHEN OTHERS;

	g_mux : mux2t1_N
	PORT MAP(
		i_S => i_En,
		i_D0 => x"00000000",
		i_D1 => decoderOut,
		o_O => o_Out);

END mixed;